* 
.subckt PM_CMOM1%P 3 4 31 32 59 60 87 88 115 116 143 144 171 172 199 200 227 228
+ 255 256 283 284 311 312 339 340 367 368 374 395 396 423 424 451 452 479 480 507
+ 508 535 536 561 563 586 612 638 664 690 716 742 768 794 820 846 872 898 924
+ 950 976 1002 1028 1054 1080 1106 1132 1158 1184 1210 1236 1262 1288 1314 1340
+ 1366 1392 1418 1444 1470 1496 1522 1548 1574 1600 VSS
c82 1600 VSS 0.00538176f
c83 1574 VSS 0.00538176f
c84 1548 VSS 0.00538176f
c85 1522 VSS 0.00538176f
c86 1496 VSS 0.00538176f
c87 1470 VSS 0.00538176f
c88 1444 VSS 0.00538176f
c89 1418 VSS 0.00538176f
c90 1392 VSS 0.00538176f
c91 1366 VSS 0.00538176f
c92 1340 VSS 0.00538176f
c93 1314 VSS 0.00538176f
c94 1288 VSS 0.00538176f
c95 1262 VSS 0.00538176f
c96 1236 VSS 0.00538176f
c97 1210 VSS 0.00538176f
c98 1184 VSS 0.00538176f
c99 1158 VSS 0.00538176f
c100 1132 VSS 0.00538176f
c101 1106 VSS 0.00538176f
c102 1080 VSS 0.226444f
c103 1054 VSS 0.226444f
c104 1028 VSS 0.226444f
c105 1002 VSS 0.226444f
c106 976 VSS 0.226444f
c107 950 VSS 0.226444f
c108 924 VSS 0.226444f
c109 898 VSS 0.226444f
c110 872 VSS 0.226444f
c111 846 VSS 0.226444f
c112 820 VSS 0.226444f
c113 794 VSS 0.226444f
c114 768 VSS 0.226444f
c115 742 VSS 0.226444f
c116 716 VSS 0.226444f
c117 690 VSS 0.226444f
c118 664 VSS 0.226444f
c119 638 VSS 0.226444f
c120 612 VSS 0.226444f
c121 586 VSS 0.226444f
c122 561 VSS 0.743111f
c123 560 VSS 0.0164286f
c124 536 VSS 0.00398955f
c125 535 VSS 0.0025948f
c126 533 VSS 0.0149296f
c127 532 VSS 0.00479925f
c128 508 VSS 0.00398955f
c129 507 VSS 0.0025948f
c130 505 VSS 0.00426556f
c131 504 VSS 0.00479925f
c132 480 VSS 0.00398955f
c133 479 VSS 0.0025948f
c134 477 VSS 0.00426556f
c135 476 VSS 0.00479925f
c136 452 VSS 0.00398955f
c137 451 VSS 0.0025948f
c138 449 VSS 0.00426556f
c139 448 VSS 0.00479925f
c140 424 VSS 0.00398955f
c141 423 VSS 0.0025948f
c142 421 VSS 0.00426556f
c143 420 VSS 0.00479925f
c144 396 VSS 0.00398955f
c145 395 VSS 0.0025948f
c146 393 VSS 0.00426556f
c147 392 VSS 0.00479925f
c148 368 VSS 0.00398955f
c149 367 VSS 0.0025948f
c150 365 VSS 0.00426556f
c151 364 VSS 0.00479925f
c152 340 VSS 0.00398955f
c153 339 VSS 0.0025948f
c154 337 VSS 0.00426556f
c155 336 VSS 0.00479925f
c156 312 VSS 0.00398955f
c157 311 VSS 0.0025948f
c158 309 VSS 0.00426556f
c159 308 VSS 0.00479925f
c160 284 VSS 0.00398955f
c161 283 VSS 0.0025948f
c162 281 VSS 0.00426556f
c163 280 VSS 0.00479925f
c164 256 VSS 0.00398955f
c165 255 VSS 0.0025948f
c166 253 VSS 0.00426556f
c167 252 VSS 0.00479925f
c168 228 VSS 0.00398955f
c169 227 VSS 0.0025948f
c170 225 VSS 0.00426556f
c171 224 VSS 0.00479925f
c172 200 VSS 0.00398955f
c173 199 VSS 0.0025948f
c174 197 VSS 0.00426556f
c175 196 VSS 0.00479925f
c176 172 VSS 0.00398955f
c177 171 VSS 0.0025948f
c178 169 VSS 0.00426556f
c179 168 VSS 0.00479925f
c180 144 VSS 0.00398955f
c181 143 VSS 0.0025948f
c182 141 VSS 0.00426556f
c183 140 VSS 0.00479925f
c184 116 VSS 0.00398955f
c185 115 VSS 0.0025948f
c186 113 VSS 0.00426556f
c187 112 VSS 0.00479925f
c188 88 VSS 0.00398955f
c189 87 VSS 0.0025948f
c190 85 VSS 0.00426556f
c191 84 VSS 0.00479925f
c192 60 VSS 0.00398955f
c193 59 VSS 0.0025948f
c194 57 VSS 0.00426556f
c195 56 VSS 0.00479925f
c196 32 VSS 0.00398955f
c197 31 VSS 0.0025948f
c198 29 VSS 0.00426556f
c199 28 VSS 0.0164286f
c200 4 VSS 0.00398955f
c201 3 VSS 0.0025948f
c202 1 VSS 0.0149296f
r203 1619 1622 0.688159
r204 1616 1619 0.688159
r205 1613 1616 0.688159
r206 1610 1613 0.688159
r207 1607 1610 0.688159
r208 1604 1607 0.682697
r209 1600 1604 0.679966
r210 1593 1596 0.688159
r211 1590 1593 0.688159
r212 1587 1590 0.688159
r213 1584 1587 0.688159
r214 1581 1584 0.688159
r215 1578 1581 0.682697
r216 1574 1578 0.679966
r217 1567 1570 0.688159
r218 1564 1567 0.688159
r219 1561 1564 0.688159
r220 1558 1561 0.688159
r221 1555 1558 0.688159
r222 1552 1555 0.682697
r223 1548 1552 0.679966
r224 1541 1544 0.688159
r225 1538 1541 0.688159
r226 1535 1538 0.688159
r227 1532 1535 0.688159
r228 1529 1532 0.688159
r229 1526 1529 0.682697
r230 1522 1526 0.679966
r231 1515 1518 0.688159
r232 1512 1515 0.688159
r233 1509 1512 0.688159
r234 1506 1509 0.688159
r235 1503 1506 0.688159
r236 1500 1503 0.682697
r237 1496 1500 0.679966
r238 1489 1492 0.688159
r239 1486 1489 0.688159
r240 1483 1486 0.688159
r241 1480 1483 0.688159
r242 1477 1480 0.688159
r243 1474 1477 0.682697
r244 1470 1474 0.679966
r245 1463 1466 0.688159
r246 1460 1463 0.688159
r247 1457 1460 0.688159
r248 1454 1457 0.688159
r249 1451 1454 0.688159
r250 1448 1451 0.682697
r251 1444 1448 0.679966
r252 1437 1440 0.688159
r253 1434 1437 0.688159
r254 1431 1434 0.688159
r255 1428 1431 0.688159
r256 1425 1428 0.688159
r257 1422 1425 0.682697
r258 1418 1422 0.679966
r259 1411 1414 0.688159
r260 1408 1411 0.688159
r261 1405 1408 0.688159
r262 1402 1405 0.688159
r263 1399 1402 0.688159
r264 1396 1399 0.682697
r265 1392 1396 0.679966
r266 1385 1388 0.688159
r267 1382 1385 0.688159
r268 1379 1382 0.688159
r269 1376 1379 0.688159
r270 1373 1376 0.688159
r271 1370 1373 0.682697
r272 1366 1370 0.679966
r273 1359 1362 0.688159
r274 1356 1359 0.688159
r275 1353 1356 0.688159
r276 1350 1353 0.688159
r277 1347 1350 0.688159
r278 1344 1347 0.682697
r279 1340 1344 0.679966
r280 1333 1336 0.688159
r281 1330 1333 0.688159
r282 1327 1330 0.688159
r283 1324 1327 0.688159
r284 1321 1324 0.688159
r285 1318 1321 0.682697
r286 1314 1318 0.679966
r287 1307 1310 0.688159
r288 1304 1307 0.688159
r289 1301 1304 0.688159
r290 1298 1301 0.688159
r291 1295 1298 0.688159
r292 1292 1295 0.682697
r293 1288 1292 0.679966
r294 1281 1284 0.688159
r295 1278 1281 0.688159
r296 1275 1278 0.688159
r297 1272 1275 0.688159
r298 1269 1272 0.688159
r299 1266 1269 0.682697
r300 1262 1266 0.679966
r301 1255 1258 0.688159
r302 1252 1255 0.688159
r303 1249 1252 0.688159
r304 1246 1249 0.688159
r305 1243 1246 0.688159
r306 1240 1243 0.682697
r307 1236 1240 0.679966
r308 1229 1232 0.688159
r309 1226 1229 0.688159
r310 1223 1226 0.688159
r311 1220 1223 0.688159
r312 1217 1220 0.688159
r313 1214 1217 0.682697
r314 1210 1214 0.679966
r315 1203 1206 0.688159
r316 1200 1203 0.688159
r317 1197 1200 0.688159
r318 1194 1197 0.688159
r319 1191 1194 0.688159
r320 1188 1191 0.682697
r321 1184 1188 0.679966
r322 1177 1180 0.688159
r323 1174 1177 0.688159
r324 1171 1174 0.688159
r325 1168 1171 0.688159
r326 1165 1168 0.688159
r327 1162 1165 0.682697
r328 1158 1162 0.679966
r329 1151 1154 0.688159
r330 1148 1151 0.688159
r331 1145 1148 0.688159
r332 1142 1145 0.688159
r333 1139 1142 0.688159
r334 1136 1139 0.682697
r335 1132 1136 0.679966
r336 1125 1128 0.688159
r337 1122 1125 0.688159
r338 1119 1122 0.688159
r339 1116 1119 0.688159
r340 1113 1116 0.688159
r341 1110 1113 0.682697
r342 1106 1110 0.679966
r343 1102 1622 2.33333
r344 1099 1102 1.13284
r345 1099 1619 2.33333
r346 1096 1099 1.13284
r347 1096 1616 2.33333
r348 1093 1096 1.13284
r349 1093 1613 2.33333
r350 1090 1093 1.13284
r351 1090 1610 2.33333
r352 1087 1090 1.13284
r353 1087 1607 2.33333
r354 1084 1087 1.12385
r355 1084 1604 2.33333
r356 1080 1084 1.11935
r357 1080 1600 2.33333
r358 1076 1596 2.33333
r359 1073 1076 1.13284
r360 1073 1593 2.33333
r361 1070 1073 1.13284
r362 1070 1590 2.33333
r363 1067 1070 1.13284
r364 1067 1587 2.33333
r365 1064 1067 1.13284
r366 1064 1584 2.33333
r367 1061 1064 1.13284
r368 1061 1581 2.33333
r369 1058 1061 1.12385
r370 1058 1578 2.33333
r371 1054 1058 1.11935
r372 1054 1574 2.33333
r373 1050 1570 2.33333
r374 1047 1050 1.13284
r375 1047 1567 2.33333
r376 1044 1047 1.13284
r377 1044 1564 2.33333
r378 1041 1044 1.13284
r379 1041 1561 2.33333
r380 1038 1041 1.13284
r381 1038 1558 2.33333
r382 1035 1038 1.13284
r383 1035 1555 2.33333
r384 1032 1035 1.12385
r385 1032 1552 2.33333
r386 1028 1032 1.11935
r387 1028 1548 2.33333
r388 1024 1544 2.33333
r389 1021 1024 1.13284
r390 1021 1541 2.33333
r391 1018 1021 1.13284
r392 1018 1538 2.33333
r393 1015 1018 1.13284
r394 1015 1535 2.33333
r395 1012 1015 1.13284
r396 1012 1532 2.33333
r397 1009 1012 1.13284
r398 1009 1529 2.33333
r399 1006 1009 1.12385
r400 1006 1526 2.33333
r401 1002 1006 1.11935
r402 1002 1522 2.33333
r403 998 1518 2.33333
r404 995 998 1.13284
r405 995 1515 2.33333
r406 992 995 1.13284
r407 992 1512 2.33333
r408 989 992 1.13284
r409 989 1509 2.33333
r410 986 989 1.13284
r411 986 1506 2.33333
r412 983 986 1.13284
r413 983 1503 2.33333
r414 980 983 1.12385
r415 980 1500 2.33333
r416 976 980 1.11935
r417 976 1496 2.33333
r418 972 1492 2.33333
r419 969 972 1.13284
r420 969 1489 2.33333
r421 966 969 1.13284
r422 966 1486 2.33333
r423 963 966 1.13284
r424 963 1483 2.33333
r425 960 963 1.13284
r426 960 1480 2.33333
r427 957 960 1.13284
r428 957 1477 2.33333
r429 954 957 1.12385
r430 954 1474 2.33333
r431 950 954 1.11935
r432 950 1470 2.33333
r433 946 1466 2.33333
r434 943 946 1.13284
r435 943 1463 2.33333
r436 940 943 1.13284
r437 940 1460 2.33333
r438 937 940 1.13284
r439 937 1457 2.33333
r440 934 937 1.13284
r441 934 1454 2.33333
r442 931 934 1.13284
r443 931 1451 2.33333
r444 928 931 1.12385
r445 928 1448 2.33333
r446 924 928 1.11935
r447 924 1444 2.33333
r448 920 1440 2.33333
r449 917 920 1.13284
r450 917 1437 2.33333
r451 914 917 1.13284
r452 914 1434 2.33333
r453 911 914 1.13284
r454 911 1431 2.33333
r455 908 911 1.13284
r456 908 1428 2.33333
r457 905 908 1.13284
r458 905 1425 2.33333
r459 902 905 1.12385
r460 902 1422 2.33333
r461 898 902 1.11935
r462 898 1418 2.33333
r463 894 1414 2.33333
r464 891 894 1.13284
r465 891 1411 2.33333
r466 888 891 1.13284
r467 888 1408 2.33333
r468 885 888 1.13284
r469 885 1405 2.33333
r470 882 885 1.13284
r471 882 1402 2.33333
r472 879 882 1.13284
r473 879 1399 2.33333
r474 876 879 1.12385
r475 876 1396 2.33333
r476 872 876 1.11935
r477 872 1392 2.33333
r478 868 1388 2.33333
r479 865 868 1.13284
r480 865 1385 2.33333
r481 862 865 1.13284
r482 862 1382 2.33333
r483 859 862 1.13284
r484 859 1379 2.33333
r485 856 859 1.13284
r486 856 1376 2.33333
r487 853 856 1.13284
r488 853 1373 2.33333
r489 850 853 1.12385
r490 850 1370 2.33333
r491 846 850 1.11935
r492 846 1366 2.33333
r493 842 1362 2.33333
r494 839 842 1.13284
r495 839 1359 2.33333
r496 836 839 1.13284
r497 836 1356 2.33333
r498 833 836 1.13284
r499 833 1353 2.33333
r500 830 833 1.13284
r501 830 1350 2.33333
r502 827 830 1.13284
r503 827 1347 2.33333
r504 824 827 1.12385
r505 824 1344 2.33333
r506 820 824 1.11935
r507 820 1340 2.33333
r508 816 1336 2.33333
r509 813 816 1.13284
r510 813 1333 2.33333
r511 810 813 1.13284
r512 810 1330 2.33333
r513 807 810 1.13284
r514 807 1327 2.33333
r515 804 807 1.13284
r516 804 1324 2.33333
r517 801 804 1.13284
r518 801 1321 2.33333
r519 798 801 1.12385
r520 798 1318 2.33333
r521 794 798 1.11935
r522 794 1314 2.33333
r523 790 1310 2.33333
r524 787 790 1.13284
r525 787 1307 2.33333
r526 784 787 1.13284
r527 784 1304 2.33333
r528 781 784 1.13284
r529 781 1301 2.33333
r530 778 781 1.13284
r531 778 1298 2.33333
r532 775 778 1.13284
r533 775 1295 2.33333
r534 772 775 1.12385
r535 772 1292 2.33333
r536 768 772 1.11935
r537 768 1288 2.33333
r538 764 1284 2.33333
r539 761 764 1.13284
r540 761 1281 2.33333
r541 758 761 1.13284
r542 758 1278 2.33333
r543 755 758 1.13284
r544 755 1275 2.33333
r545 752 755 1.13284
r546 752 1272 2.33333
r547 749 752 1.13284
r548 749 1269 2.33333
r549 746 749 1.12385
r550 746 1266 2.33333
r551 742 746 1.11935
r552 742 1262 2.33333
r553 738 1258 2.33333
r554 735 738 1.13284
r555 735 1255 2.33333
r556 732 735 1.13284
r557 732 1252 2.33333
r558 729 732 1.13284
r559 729 1249 2.33333
r560 726 729 1.13284
r561 726 1246 2.33333
r562 723 726 1.13284
r563 723 1243 2.33333
r564 720 723 1.12385
r565 720 1240 2.33333
r566 716 720 1.11935
r567 716 1236 2.33333
r568 712 1232 2.33333
r569 709 712 1.13284
r570 709 1229 2.33333
r571 706 709 1.13284
r572 706 1226 2.33333
r573 703 706 1.13284
r574 703 1223 2.33333
r575 700 703 1.13284
r576 700 1220 2.33333
r577 697 700 1.13284
r578 697 1217 2.33333
r579 694 697 1.12385
r580 694 1214 2.33333
r581 690 694 1.11935
r582 690 1210 2.33333
r583 686 1206 2.33333
r584 683 686 1.13284
r585 683 1203 2.33333
r586 680 683 1.13284
r587 680 1200 2.33333
r588 677 680 1.13284
r589 677 1197 2.33333
r590 674 677 1.13284
r591 674 1194 2.33333
r592 671 674 1.13284
r593 671 1191 2.33333
r594 668 671 1.12385
r595 668 1188 2.33333
r596 664 668 1.11935
r597 664 1184 2.33333
r598 660 1180 2.33333
r599 657 660 1.13284
r600 657 1177 2.33333
r601 654 657 1.13284
r602 654 1174 2.33333
r603 651 654 1.13284
r604 651 1171 2.33333
r605 648 651 1.13284
r606 648 1168 2.33333
r607 645 648 1.13284
r608 645 1165 2.33333
r609 642 645 1.12385
r610 642 1162 2.33333
r611 638 642 1.11935
r612 638 1158 2.33333
r613 634 1154 2.33333
r614 631 634 1.13284
r615 631 1151 2.33333
r616 628 631 1.13284
r617 628 1148 2.33333
r618 625 628 1.13284
r619 625 1145 2.33333
r620 622 625 1.13284
r621 622 1142 2.33333
r622 619 622 1.13284
r623 619 1139 2.33333
r624 616 619 1.12385
r625 616 1136 2.33333
r626 612 616 1.11935
r627 612 1132 2.33333
r628 608 1128 2.33333
r629 605 608 1.13284
r630 605 1125 2.33333
r631 602 605 1.13284
r632 602 1122 2.33333
r633 599 602 1.13284
r634 599 1119 2.33333
r635 596 599 1.13284
r636 596 1116 2.33333
r637 593 596 1.13284
r638 593 1113 2.33333
r639 590 593 1.12385
r640 590 1110 2.33333
r641 586 590 1.11935
r642 586 1106 2.33333
r643 583 584 0.0895699
r644 582 583 0.0895699
r645 581 582 0.0895699
r646 580 581 0.0895699
r647 579 580 0.0895699
r648 578 579 0.0895699
r649 577 578 0.0895699
r650 576 577 0.0895699
r651 575 576 0.0895699
r652 574 575 0.0895699
r653 573 574 0.0895699
r654 572 573 0.0895699
r655 571 572 0.0895699
r656 570 571 0.0895699
r657 569 570 0.0895699
r658 568 569 0.0895699
r659 567 568 0.0895699
r660 566 567 0.0895699
r661 565 566 0.0895699
r662 563 565 0.0557081
r663 561 584 0.0229386
r664 559 560 0.273079
r665 558 1622 2.33333
r666 557 559 0.330425
r667 557 558 2.33333
r668 555 558 0.688159
r669 555 1619 2.33333
r670 554 557 0.688159
r671 554 555 2.33333
r672 552 555 0.688159
r673 552 1616 2.33333
r674 551 554 0.688159
r675 551 552 2.33333
r676 549 552 0.688159
r677 549 1613 2.33333
r678 548 551 0.688159
r679 548 549 2.33333
r680 546 549 0.688159
r681 546 1610 2.33333
r682 545 548 0.688159
r683 545 546 2.33333
r684 543 546 0.688159
r685 543 1607 2.33333
r686 542 545 0.688159
r687 542 543 2.33333
r688 540 543 0.682697
r689 540 1604 2.33333
r690 539 542 0.682697
r691 539 540 2.33333
r692 536 540 0.679966
r693 536 1600 2.33333
r694 535 539 0.679966
r695 535 536 2.33333
r696 533 584 0.0950558
r697 533 560 0.273079
r698 531 532 0.273079
r699 530 1596 2.33333
r700 529 531 0.330425
r701 529 530 2.33333
r702 527 530 0.688159
r703 527 1593 2.33333
r704 526 529 0.688159
r705 526 527 2.33333
r706 524 527 0.688159
r707 524 1590 2.33333
r708 523 526 0.688159
r709 523 524 2.33333
r710 521 524 0.688159
r711 521 1587 2.33333
r712 520 523 0.688159
r713 520 521 2.33333
r714 518 521 0.688159
r715 518 1584 2.33333
r716 517 520 0.688159
r717 517 518 2.33333
r718 515 518 0.688159
r719 515 1581 2.33333
r720 514 517 0.688159
r721 514 515 2.33333
r722 512 515 0.682697
r723 512 1578 2.33333
r724 511 514 0.682697
r725 511 512 2.33333
r726 508 512 0.679966
r727 508 1574 2.33333
r728 507 511 0.679966
r729 507 508 2.33333
r730 505 583 0.0950558
r731 505 532 0.273079
r732 503 504 0.273079
r733 502 1570 2.33333
r734 501 503 0.330425
r735 501 502 2.33333
r736 499 502 0.688159
r737 499 1567 2.33333
r738 498 501 0.688159
r739 498 499 2.33333
r740 496 499 0.688159
r741 496 1564 2.33333
r742 495 498 0.688159
r743 495 496 2.33333
r744 493 496 0.688159
r745 493 1561 2.33333
r746 492 495 0.688159
r747 492 493 2.33333
r748 490 493 0.688159
r749 490 1558 2.33333
r750 489 492 0.688159
r751 489 490 2.33333
r752 487 490 0.688159
r753 487 1555 2.33333
r754 486 489 0.688159
r755 486 487 2.33333
r756 484 487 0.682697
r757 484 1552 2.33333
r758 483 486 0.682697
r759 483 484 2.33333
r760 480 484 0.679966
r761 480 1548 2.33333
r762 479 483 0.679966
r763 479 480 2.33333
r764 477 582 0.0950558
r765 477 504 0.273079
r766 475 476 0.273079
r767 474 1544 2.33333
r768 473 475 0.330425
r769 473 474 2.33333
r770 471 474 0.688159
r771 471 1541 2.33333
r772 470 473 0.688159
r773 470 471 2.33333
r774 468 471 0.688159
r775 468 1538 2.33333
r776 467 470 0.688159
r777 467 468 2.33333
r778 465 468 0.688159
r779 465 1535 2.33333
r780 464 467 0.688159
r781 464 465 2.33333
r782 462 465 0.688159
r783 462 1532 2.33333
r784 461 464 0.688159
r785 461 462 2.33333
r786 459 462 0.688159
r787 459 1529 2.33333
r788 458 461 0.688159
r789 458 459 2.33333
r790 456 459 0.682697
r791 456 1526 2.33333
r792 455 458 0.682697
r793 455 456 2.33333
r794 452 456 0.679966
r795 452 1522 2.33333
r796 451 455 0.679966
r797 451 452 2.33333
r798 449 581 0.0950558
r799 449 476 0.273079
r800 447 448 0.273079
r801 446 1518 2.33333
r802 445 447 0.330425
r803 445 446 2.33333
r804 443 446 0.688159
r805 443 1515 2.33333
r806 442 445 0.688159
r807 442 443 2.33333
r808 440 443 0.688159
r809 440 1512 2.33333
r810 439 442 0.688159
r811 439 440 2.33333
r812 437 440 0.688159
r813 437 1509 2.33333
r814 436 439 0.688159
r815 436 437 2.33333
r816 434 437 0.688159
r817 434 1506 2.33333
r818 433 436 0.688159
r819 433 434 2.33333
r820 431 434 0.688159
r821 431 1503 2.33333
r822 430 433 0.688159
r823 430 431 2.33333
r824 428 431 0.682697
r825 428 1500 2.33333
r826 427 430 0.682697
r827 427 428 2.33333
r828 424 428 0.679966
r829 424 1496 2.33333
r830 423 427 0.679966
r831 423 424 2.33333
r832 421 580 0.0950558
r833 421 448 0.273079
r834 419 420 0.273079
r835 418 1492 2.33333
r836 417 419 0.330425
r837 417 418 2.33333
r838 415 418 0.688159
r839 415 1489 2.33333
r840 414 417 0.688159
r841 414 415 2.33333
r842 412 415 0.688159
r843 412 1486 2.33333
r844 411 414 0.688159
r845 411 412 2.33333
r846 409 412 0.688159
r847 409 1483 2.33333
r848 408 411 0.688159
r849 408 409 2.33333
r850 406 409 0.688159
r851 406 1480 2.33333
r852 405 408 0.688159
r853 405 406 2.33333
r854 403 406 0.688159
r855 403 1477 2.33333
r856 402 405 0.688159
r857 402 403 2.33333
r858 400 403 0.682697
r859 400 1474 2.33333
r860 399 402 0.682697
r861 399 400 2.33333
r862 396 400 0.679966
r863 396 1470 2.33333
r864 395 399 0.679966
r865 395 396 2.33333
r866 393 579 0.0950558
r867 393 420 0.273079
r868 391 392 0.273079
r869 390 1466 2.33333
r870 389 391 0.330425
r871 389 390 2.33333
r872 387 390 0.688159
r873 387 1463 2.33333
r874 386 389 0.688159
r875 386 387 2.33333
r876 384 387 0.688159
r877 384 1460 2.33333
r878 383 386 0.688159
r879 383 384 2.33333
r880 381 384 0.688159
r881 381 1457 2.33333
r882 380 383 0.688159
r883 380 381 2.33333
r884 378 381 0.688159
r885 378 1454 2.33333
r886 377 380 0.688159
r887 377 378 2.33333
r888 375 378 0.688159
r889 375 1451 2.33333
r890 374 377 0.688159
r891 374 375 2.33333
r892 372 375 0.682697
r893 372 1448 2.33333
r894 371 374 0.682697
r895 371 372 2.33333
r896 368 372 0.679966
r897 368 1444 2.33333
r898 367 371 0.679966
r899 367 368 2.33333
r900 365 578 0.0950558
r901 365 392 0.273079
r902 363 364 0.273079
r903 362 1440 2.33333
r904 361 363 0.330425
r905 361 362 2.33333
r906 359 362 0.688159
r907 359 1437 2.33333
r908 358 361 0.688159
r909 358 359 2.33333
r910 356 359 0.688159
r911 356 1434 2.33333
r912 355 358 0.688159
r913 355 356 2.33333
r914 353 356 0.688159
r915 353 1431 2.33333
r916 352 355 0.688159
r917 352 353 2.33333
r918 350 353 0.688159
r919 350 1428 2.33333
r920 349 352 0.688159
r921 349 350 2.33333
r922 347 350 0.688159
r923 347 1425 2.33333
r924 346 349 0.688159
r925 346 347 2.33333
r926 344 347 0.682697
r927 344 1422 2.33333
r928 343 346 0.682697
r929 343 344 2.33333
r930 340 344 0.679966
r931 340 1418 2.33333
r932 339 343 0.679966
r933 339 340 2.33333
r934 337 577 0.0950558
r935 337 364 0.273079
r936 335 336 0.273079
r937 334 1414 2.33333
r938 333 335 0.330425
r939 333 334 2.33333
r940 331 334 0.688159
r941 331 1411 2.33333
r942 330 333 0.688159
r943 330 331 2.33333
r944 328 331 0.688159
r945 328 1408 2.33333
r946 327 330 0.688159
r947 327 328 2.33333
r948 325 328 0.688159
r949 325 1405 2.33333
r950 324 327 0.688159
r951 324 325 2.33333
r952 322 325 0.688159
r953 322 1402 2.33333
r954 321 324 0.688159
r955 321 322 2.33333
r956 319 322 0.688159
r957 319 1399 2.33333
r958 318 321 0.688159
r959 318 319 2.33333
r960 316 319 0.682697
r961 316 1396 2.33333
r962 315 318 0.682697
r963 315 316 2.33333
r964 312 316 0.679966
r965 312 1392 2.33333
r966 311 315 0.679966
r967 311 312 2.33333
r968 309 576 0.0950558
r969 309 336 0.273079
r970 307 308 0.273079
r971 306 1388 2.33333
r972 305 307 0.330425
r973 305 306 2.33333
r974 303 306 0.688159
r975 303 1385 2.33333
r976 302 305 0.688159
r977 302 303 2.33333
r978 300 303 0.688159
r979 300 1382 2.33333
r980 299 302 0.688159
r981 299 300 2.33333
r982 297 300 0.688159
r983 297 1379 2.33333
r984 296 299 0.688159
r985 296 297 2.33333
r986 294 297 0.688159
r987 294 1376 2.33333
r988 293 296 0.688159
r989 293 294 2.33333
r990 291 294 0.688159
r991 291 1373 2.33333
r992 290 293 0.688159
r993 290 291 2.33333
r994 288 291 0.682697
r995 288 1370 2.33333
r996 287 290 0.682697
r997 287 288 2.33333
r998 284 288 0.679966
r999 284 1366 2.33333
r1000 283 287 0.679966
r1001 283 284 2.33333
r1002 281 575 0.0950558
r1003 281 308 0.273079
r1004 279 280 0.273079
r1005 278 1362 2.33333
r1006 277 279 0.330425
r1007 277 278 2.33333
r1008 275 278 0.688159
r1009 275 1359 2.33333
r1010 274 277 0.688159
r1011 274 275 2.33333
r1012 272 275 0.688159
r1013 272 1356 2.33333
r1014 271 274 0.688159
r1015 271 272 2.33333
r1016 269 272 0.688159
r1017 269 1353 2.33333
r1018 268 271 0.688159
r1019 268 269 2.33333
r1020 266 269 0.688159
r1021 266 1350 2.33333
r1022 265 268 0.688159
r1023 265 266 2.33333
r1024 263 266 0.688159
r1025 263 1347 2.33333
r1026 262 265 0.688159
r1027 262 263 2.33333
r1028 260 263 0.682697
r1029 260 1344 2.33333
r1030 259 262 0.682697
r1031 259 260 2.33333
r1032 256 260 0.679966
r1033 256 1340 2.33333
r1034 255 259 0.679966
r1035 255 256 2.33333
r1036 253 574 0.0950558
r1037 253 280 0.273079
r1038 251 252 0.273079
r1039 250 1336 2.33333
r1040 249 251 0.330425
r1041 249 250 2.33333
r1042 247 250 0.688159
r1043 247 1333 2.33333
r1044 246 249 0.688159
r1045 246 247 2.33333
r1046 244 247 0.688159
r1047 244 1330 2.33333
r1048 243 246 0.688159
r1049 243 244 2.33333
r1050 241 244 0.688159
r1051 241 1327 2.33333
r1052 240 243 0.688159
r1053 240 241 2.33333
r1054 238 241 0.688159
r1055 238 1324 2.33333
r1056 237 240 0.688159
r1057 237 238 2.33333
r1058 235 238 0.688159
r1059 235 1321 2.33333
r1060 234 237 0.688159
r1061 234 235 2.33333
r1062 232 235 0.682697
r1063 232 1318 2.33333
r1064 231 234 0.682697
r1065 231 232 2.33333
r1066 228 232 0.679966
r1067 228 1314 2.33333
r1068 227 231 0.679966
r1069 227 228 2.33333
r1070 225 573 0.0950558
r1071 225 252 0.273079
r1072 223 224 0.273079
r1073 222 1310 2.33333
r1074 221 223 0.330425
r1075 221 222 2.33333
r1076 219 222 0.688159
r1077 219 1307 2.33333
r1078 218 221 0.688159
r1079 218 219 2.33333
r1080 216 219 0.688159
r1081 216 1304 2.33333
r1082 215 218 0.688159
r1083 215 216 2.33333
r1084 213 216 0.688159
r1085 213 1301 2.33333
r1086 212 215 0.688159
r1087 212 213 2.33333
r1088 210 213 0.688159
r1089 210 1298 2.33333
r1090 209 212 0.688159
r1091 209 210 2.33333
r1092 207 210 0.688159
r1093 207 1295 2.33333
r1094 206 209 0.688159
r1095 206 207 2.33333
r1096 204 207 0.682697
r1097 204 1292 2.33333
r1098 203 206 0.682697
r1099 203 204 2.33333
r1100 200 204 0.679966
r1101 200 1288 2.33333
r1102 199 203 0.679966
r1103 199 200 2.33333
r1104 197 572 0.0950558
r1105 197 224 0.273079
r1106 195 196 0.273079
r1107 194 1284 2.33333
r1108 193 195 0.330425
r1109 193 194 2.33333
r1110 191 194 0.688159
r1111 191 1281 2.33333
r1112 190 193 0.688159
r1113 190 191 2.33333
r1114 188 191 0.688159
r1115 188 1278 2.33333
r1116 187 190 0.688159
r1117 187 188 2.33333
r1118 185 188 0.688159
r1119 185 1275 2.33333
r1120 184 187 0.688159
r1121 184 185 2.33333
r1122 182 185 0.688159
r1123 182 1272 2.33333
r1124 181 184 0.688159
r1125 181 182 2.33333
r1126 179 182 0.688159
r1127 179 1269 2.33333
r1128 178 181 0.688159
r1129 178 179 2.33333
r1130 176 179 0.682697
r1131 176 1266 2.33333
r1132 175 178 0.682697
r1133 175 176 2.33333
r1134 172 176 0.679966
r1135 172 1262 2.33333
r1136 171 175 0.679966
r1137 171 172 2.33333
r1138 169 571 0.0950558
r1139 169 196 0.273079
r1140 167 168 0.273079
r1141 166 1258 2.33333
r1142 165 167 0.330425
r1143 165 166 2.33333
r1144 163 166 0.688159
r1145 163 1255 2.33333
r1146 162 165 0.688159
r1147 162 163 2.33333
r1148 160 163 0.688159
r1149 160 1252 2.33333
r1150 159 162 0.688159
r1151 159 160 2.33333
r1152 157 160 0.688159
r1153 157 1249 2.33333
r1154 156 159 0.688159
r1155 156 157 2.33333
r1156 52 157 0.688159
r1157 154 1246 2.33333
r1158 153 156 0.688159
r1159 153 154 2.33333
r1160 151 154 0.688159
r1161 151 1243 2.33333
r1162 150 153 0.688159
r1163 150 151 2.33333
r1164 148 151 0.682697
r1165 148 1240 2.33333
r1166 147 150 0.682697
r1167 147 148 2.33333
r1168 144 148 0.679966
r1169 144 1236 2.33333
r1170 143 147 0.679966
r1171 143 144 2.33333
r1172 141 570 0.0950558
r1173 141 168 0.273079
r1174 139 140 0.273079
r1175 138 1232 2.33333
r1176 137 139 0.330425
r1177 137 138 2.33333
r1178 135 138 0.688159
r1179 135 1229 2.33333
r1180 134 137 0.688159
r1181 134 135 2.33333
r1182 132 135 0.688159
r1183 132 1226 2.33333
r1184 131 134 0.688159
r1185 131 132 2.33333
r1186 129 132 0.688159
r1187 129 1223 2.33333
r1188 128 131 0.688159
r1189 128 129 2.33333
r1190 126 129 0.688159
r1191 126 1220 2.33333
r1192 125 128 0.688159
r1193 125 126 2.33333
r1194 123 126 0.688159
r1195 123 1217 2.33333
r1196 122 125 0.688159
r1197 122 123 2.33333
r1198 120 123 0.682697
r1199 120 1214 2.33333
r1200 119 122 0.682697
r1201 119 120 2.33333
r1202 116 120 0.679966
r1203 116 1210 2.33333
r1204 115 119 0.679966
r1205 115 116 2.33333
r1206 113 569 0.0950558
r1207 113 140 0.273079
r1208 111 112 0.273079
r1209 110 1206 2.33333
r1210 109 111 0.330425
r1211 109 110 2.33333
r1212 107 110 0.688159
r1213 107 1203 2.33333
r1214 106 109 0.688159
r1215 106 107 2.33333
r1216 104 107 0.688159
r1217 104 1200 2.33333
r1218 103 106 0.688159
r1219 103 104 2.33333
r1220 101 104 0.688159
r1221 101 1197 2.33333
r1222 100 103 0.688159
r1223 100 101 2.33333
r1224 98 101 0.688159
r1225 98 1194 2.33333
r1226 97 100 0.688159
r1227 97 98 2.33333
r1228 95 98 0.688159
r1229 95 1191 2.33333
r1230 94 97 0.688159
r1231 94 95 2.33333
r1232 92 95 0.682697
r1233 92 1188 2.33333
r1234 91 94 0.682697
r1235 91 92 2.33333
r1236 88 92 0.679966
r1237 88 1184 2.33333
r1239 87 88 2.33333
r1240 85 568 0.0950558
r1241 85 112 0.273079
r1242 83 84 0.273079
r1243 82 1180 2.33333
r1244 81 83 0.330425
r1245 81 82 2.33333
r1246 79 82 0.688159
r1247 79 1177 2.33333
r1248 78 81 0.688159
r1249 78 79 2.33333
r1250 76 79 0.688159
r1251 76 1174 2.33333
r1252 75 78 0.688159
r1253 75 76 2.33333
r1254 73 76 0.688159
r1255 73 1171 2.33333
r1256 72 75 0.688159
r1257 72 73 2.33333
r1258 70 73 0.688159
r1259 70 1168 2.33333
r1260 69 72 0.688159
r1261 69 70 2.33333
r1262 67 70 0.688159
r1263 67 1165 2.33333
r1264 66 69 0.688159
r1265 66 67 2.33333
r1266 64 67 0.682697
r1267 64 1162 2.33333
r1268 63 66 0.682697
r1269 63 64 2.33333
r1270 60 64 0.679966
r1271 60 1158 2.33333
r1272 59 63 0.679966
r1273 59 60 2.33333
r1274 57 567 0.0950558
r1275 57 84 0.273079
r1276 55 56 0.273079
r1277 54 1154 2.33333
r1279 53 54 2.33333
r1280 51 54 0.688159
r1281 51 1151 2.33333
r1282 50 53 0.688159
r1283 50 51 2.33333
r1284 48 51 0.688159
r1285 48 1148 2.33333
r1286 47 50 0.688159
r1287 47 48 2.33333
r1288 45 48 0.688159
r1289 45 1145 2.33333
r1290 44 47 0.688159
r1291 44 45 2.33333
r1292 42 45 0.688159
r1293 42 1142 2.33333
r1294 41 44 0.688159
r1295 41 42 2.33333
r1296 39 42 0.688159
r1297 39 1139 2.33333
r1298 38 41 0.688159
r1299 38 39 2.33333
r1300 36 39 0.682697
r1301 36 1136 2.33333
r1302 35 38 0.682697
r1303 35 36 2.33333
r1304 32 36 0.679966
r1305 32 1132 2.33333
r1306 31 35 0.679966
r1307 31 32 2.33333
r1308 29 566 0.0950558
r1309 29 56 0.273079
r1310 27 28 0.273079
r1311 26 1128 2.33333
r1312 25 27 0.330425
r1313 25 26 2.33333
r1314 23 26 0.688159
r1315 23 1125 2.33333
r1316 22 25 0.688159
r1317 22 23 2.33333
r1318 20 23 0.688159
r1319 20 1122 2.33333
r1320 19 22 0.688159
r1321 19 20 2.33333
r1322 17 20 0.688159
r1323 17 1119 2.33333
r1324 16 19 0.688159
r1325 16 17 2.33333
r1326 14 17 0.688159
r1327 14 1116 2.33333
r1328 13 16 0.688159
r1329 13 14 2.33333
r1330 11 14 0.688159
r1331 11 1113 2.33333
r1332 10 13 0.688159
r1333 10 11 2.33333
r1334 8 11 0.682697
r1335 8 1110 2.33333
r1336 7 10 0.682697
r1337 7 8 2.33333
r1338 4 8 0.679966
r1339 4 1106 2.33333
r1340 3 7 0.679966
r1341 3 4 2.33333
r1342 1 565 0.0950558
r1343 1 28 0.273079
r1344 1 374 2.75698
r1345 12 6 1.7896
r1346 6 2 5.8794
r1347 2 12 3.5574
.ends



 
x_PM_CMOM1%P N_P_c_1_p N_P_c_2_p N_P_c_3_p N_P_c_4_p N_P_c_5_p N_P_c_6_p
+ N_P_c_7_p N_P_c_8_p N_P_c_9_p N_P_c_10_p N_P_c_11_p N_P_c_12_p N_P_c_13_p
+ N_P_c_14_p N_P_c_15_p N_P_c_16_p N_P_c_17_p N_P_c_18_p N_P_c_19_p N_P_c_20_p
+ N_P_c_21_p N_P_c_22_p N_P_c_23_p N_P_c_24_p N_P_c_25_p N_P_c_26_p N_P_c_27_p
+ N_P_c_28_p N_P_c_29_p N_P_c_30_p N_P_c_31_p N_P_c_32_p N_P_c_33_p N_P_c_34_p
+ N_P_c_35_p N_P_c_36_p N_P_c_37_p N_P_c_38_p N_P_c_39_p N_P_c_40_p N_P_X0_POS P
+ N_P_c_42_p N_P_c_43_p N_P_c_44_p N_P_c_45_p N_P_c_46_p N_P_c_47_p N_P_c_48_p
+ N_P_c_49_p N_P_c_50_p N_P_c_51_p N_P_c_52_p N_P_c_53_p N_P_c_54_p N_P_c_55_p
+ N_P_c_56_p N_P_c_57_p N_P_c_58_p N_P_c_59_p N_P_c_60_p N_P_c_61_p N_P_c_62_p
+ N_P_c_63_p N_P_c_64_p N_P_c_65_p N_P_c_66_p N_P_c_67_p N_P_c_68_p N_P_c_69_p
+ N_P_c_70_p N_P_c_71_p N_P_c_72_p N_P_c_73_p N_P_c_74_p N_P_c_75_p N_P_c_76_p
+ N_P_c_77_p N_P_c_78_p N_P_c_79_p N_P_c_80_p N_P_c_81_p VSS PM_CMOM1%P
cc_1 N_P_c_1_p N 2.30605f
cc_2 N_P_c_2_p N 3.27983f
cc_3 N_P_c_3_p N 2.2952f
cc_4 N_P_c_4_p N 3.28318f
cc_5 N_P_c_5_p N 2.2952f
cc_6 N_P_c_6_p N 3.28318f
cc_7 N_P_c_7_p N 2.2952f
cc_8 N_P_c_8_p N 3.28318f
cc_9 N_P_c_9_p N 2.2952f
cc_10 N_P_c_10_p N 3.28318f
cc_11 N_P_c_11_p N 2.2952f
cc_12 N_P_c_12_p N 3.28318f
cc_13 N_P_c_13_p N 2.2952f
cc_14 N_P_c_14_p N 3.28318f
cc_15 N_P_c_15_p N 2.2952f
cc_16 N_P_c_16_p N 3.28318f
cc_17 N_P_c_17_p N 2.2952f
cc_18 N_P_c_18_p N 3.28318f
cc_19 N_P_c_19_p N 2.2952f
cc_20 N_P_c_20_p N 3.28318f
cc_21 N_P_c_21_p N 2.2952f
cc_22 N_P_c_22_p N 3.28318f
cc_23 N_P_c_23_p N 2.2952f
cc_24 N_P_c_24_p N 3.28318f
cc_25 N_P_c_25_p N 2.2952f
cc_26 N_P_c_26_p N 3.28318f
cc_27 N_P_c_27_p N 2.2952f
cc_28 N_P_c_28_p N 3.28318f
cc_29 N_P_c_29_p N 2.2952f
cc_30 N_P_c_30_p N 3.28318f
cc_31 N_P_c_31_p N 2.2952f
cc_32 N_P_c_32_p N 3.28318f
cc_33 N_P_c_33_p N 2.2952f
cc_34 N_P_c_34_p N 3.28318f
cc_35 N_P_c_35_p N 2.2952f
cc_36 N_P_c_36_p N 3.28318f
cc_37 N_P_c_37_p N 2.2952f
cc_38 N_P_c_38_p N 3.28318f
cc_39 N_P_c_39_p N 2.30605f
cc_40 N_P_c_40_p N 3.27983f
cc_41 N_P_X0_POS N 0.197462f
cc_42 N_P_c_42_p N 2.95243f
cc_43 N_P_c_43_p N 2.94976f
cc_44 N_P_c_44_p N 2.94976f
cc_45 N_P_c_45_p N 2.94976f
cc_46 N_P_c_46_p N 2.94976f
cc_47 N_P_c_47_p N 2.94976f
cc_48 N_P_c_48_p N 2.94976f
cc_49 N_P_c_49_p N 2.94976f
cc_50 N_P_c_50_p N 2.94976f
cc_51 N_P_c_51_p N 2.94976f
cc_52 N_P_c_52_p N 2.94976f
cc_53 N_P_c_53_p N 2.94976f
cc_54 N_P_c_54_p N 2.94976f
cc_55 N_P_c_55_p N 2.94976f
cc_56 N_P_c_56_p N 2.94976f
cc_57 N_P_c_57_p N 2.94976f
cc_58 N_P_c_58_p N 2.94976f
cc_59 N_P_c_59_p N 2.94976f
cc_60 N_P_c_60_p N 2.94976f
cc_61 N_P_c_61_p N 2.95243f
cc_62 N_P_c_62_p N 3.2564f
cc_63 N_P_c_63_p N 3.26013f
cc_64 N_P_c_64_p N 3.26013f
cc_65 N_P_c_65_p N 3.26013f
cc_66 N_P_c_66_p N 3.26013f
cc_67 N_P_c_67_p N 3.26013f
cc_68 N_P_c_68_p N 3.26013f
cc_69 N_P_c_69_p N 3.26013f
cc_70 N_P_c_70_p N 3.26013f
cc_71 N_P_c_71_p N 3.26013f
cc_72 N_P_c_72_p N 3.26013f
cc_73 N_P_c_73_p N 3.26013f
cc_74 N_P_c_74_p N 3.26013f
cc_75 N_P_c_75_p N 3.26013f
cc_76 N_P_c_76_p N 3.26013f
cc_77 N_P_c_77_p N 3.26013f
cc_78 N_P_c_78_p N 3.26013f
cc_79 N_P_c_79_p N 3.26013f
cc_80 N_P_c_80_p N 3.26013f
cc_81 N_P_c_81_p N 3.2564f
cc_82 N_P_X0_POS 3 0.122474f
cc_83 N 3 0.00648268f
cc_84 N 52 3.26013f



